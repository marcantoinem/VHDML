library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity vhdml_top is
    port(
        clk      : in std_logic
    );
end;

architecture rtl of vhdml_top is
begin
        
end rtl;